/*******************************************************
*  AN7   AN6   AN5   AN4  | AN3   AN2   AN1   AN0
*   |     |     |     |   |  |     |     |     |
*   __    __    __    __  |  __    __    __    __
*  |__|  |__|  |__|  |__| | |__|  |__|  |__|  |__|
*  |__|. |__|. |__|. |__|.| |__|. |__|. |__|. |__|.
*      
*  | |   | |   | |   | |  |  | |   | |   | |   | |
* CA CB CC CD CE CF CG DP | CA CB CC CD CE CF CG DP
********************************************************/

/********************************************************
*              _____
*          ___|  A  |___
*         |   |-----|   |
*         | F |     | B |
*         |___|-----|___|
*          ___|  G  |___
*         |   |-----|   |
*         | E |     | C |
*         |___|_____|___|     ---
*             |  D  |        | P |
*              -----          ---
*********************************************************/

/*********************************************************
*   0     1     2     3     4     5     6     7      8     9
*   |     |     |     |     |     |     |     |      |     |  
*   __          __    __           __    __    __    __    __  
*  |  |     |   __|   __|   |__|  |__   |__      |  |__|  |__|  
*  |__|     |  |__    __|      |   __|  |__|     |  |__|   __|
*********************************************************/
module BCD_to_Cathodes (
    input [3:0] digit,
    output reg [7:0] cathode
);

  always @(digit) begin
    case (digit)
      /* dec digit      |P|G|F|E|D|C|B|A|  */
      4'd0: cathode = 8'b1_1_0_0_0_0_0_0;
      4'd1: cathode = 8'b1_1_1_1_1_0_0_1;
      4'd2: cathode = 8'b1_0_1_0_0_1_0_0;
      4'd3: cathode = 8'b1_0_1_1_0_0_0_0;
      4'd4: cathode = 8'b1_0_0_1_1_0_0_1;
      4'd5: cathode = 8'b1_0_0_1_0_0_1_0;
      4'd6: cathode = 8'b1_0_0_0_0_0_1_0;
      4'd7: cathode = 8'b1_1_1_1_1_0_0_0;
      4'd8: cathode = 8'b1_0_0_0_0_0_0_0;
      4'd9: cathode = 8'b1_0_0_1_0_0_0_0;
      /* dec digit       |P|G|F|E|D|C|B|A|  */
      4'd10: cathode = 8'b1_0_0_0_1_0_0_0; //A
      4'd11: cathode = 8'b1_0_0_0_0_0_1_1; //B
      4'd12: cathode = 8'b1_1_0_0_0_1_1_0; //C
      4'd13: cathode = 8'b1_0_1_0_0_0_0_1; //D
      4'd14: cathode = 8'b1_0_0_0_0_1_1_0; //E
      4'd15: cathode = 8'b1_0_0_0_1_1_1_0; //F
      default: cathode = 8'b1_1_1_1_1_1_1_1;
    endcase
  end


endmodule
